`ifndef DEFAULT_ENV_PKG_SVH
`define DEFAULT_ENV_PKG_SVH

  `include "default_env_config.sv"
  `include "default_env.sv"

`endif
