`ifndef DEFAULT_DEFINES_SVH
`define DEFAULT_DEFINES_SVH

`endif
