`ifndef DEFAULT_MASTER_PKG_SVH
`define DEFAULT_MASTER_PKG_SVH

  `include "default_master_config.sv"
  `include "default_master_item.sv"
  `include "default_master_sequence_lib.sv"
  `include "default_master_callbacks.sv"
  `include "default_master_sequencer.sv"
  `include "default_master_driver.sv"
  `include "default_master_monitor.sv"
  `include "default_master_analyzer.sv"
  `include "default_master_collector.sv"
  `include "default_master_adapter.sv"
  `include "default_master_agent.sv"

`endif
