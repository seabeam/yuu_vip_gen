`ifndef DEFAULT_TYPE_SV
`define DEFAULT_TYPE_SV

`endif
