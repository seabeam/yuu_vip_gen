`ifndef DEFAULT_TYPE_SVH
`define DEFAULT_TYPE_SVH

`endif
