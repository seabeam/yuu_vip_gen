`ifndef DEFAULT_SLAVE_PKG_SVH
`define DEFAULT_SLAVE_PKG_SVH

  `include "default_slave_config.sv"
  `include "default_slave_item.sv"
  `include "default_slave_sequence_lib.sv"
  `include "default_slave_callbacks.sv"
  `include "default_slave_sequencer.sv"
  `include "default_slave_driver.sv"
  `include "default_slave_monitor.sv"
  `include "default_slave_analyzer.sv"
  `include "default_slave_collector.sv"
  `include "default_slave_agent.sv"

`endif
