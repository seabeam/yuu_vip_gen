`ifndef DEFAULT_COMMON_PKG_SVH
`define DEFAULT_COMMON_PKG_SVH

  `include "default_type.sv"
  `include "default_common_agent_config.sv"
  `include "default_common_item.sv"

`endif
